<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<Root>
	<creator type="key">ConfigurationDesk 6.7</creator>
	<application>
		<Name type="key">Furuta_Acados.CDL</Name>
		<DisplayName type="key">Furuta_Acados</DisplayName>
		<Path type="key">.\Furuta_Acados</Path>
		<Component type="key">ProjectApplication</Component>
		<Type type="key">14</Type>
		<ApplicationType type="key">3</ApplicationType>
		<Flags type="key">41216</Flags>
		<ItemInfoDate type="key">28.03.2024 10:08:04</ItemInfoDate>
		<ItemInfoPath type="key">$FPATH$</ItemInfoPath>
		<ItemInfoDocs type="key"/>
		<ItemInfoDescr type="key"/>
		<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
		<Log type="key"/>
		<AddInfoDb type="key"/>
		<DatabaseID type="key">-1</DatabaseID>
		<EntityID type="key">{38C4195B-25BC-4F9C-9BEE-C705C57F89FE}</EntityID>
		<item>
			<Name type="key">WindowConfiguration.xml</Name>
			<DisplayName type="key">WindowConfiguration.xml</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">4</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{2E4118A6-4744-4C8D-913D-A2BA5616EB7F}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Device Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">33</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{9FA036FD-944E-4D16-B830-FFF1CB8C604D}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Hardware Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">19</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{CA556850-A45D-4CD2-9295-C3B4A5C94AF8}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Model Topology</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">31</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key">Model location:
C:\Users\Administrator\Furuta\Furuta_Model.slx
</Log>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{1C7AD77F-05D3-4ECB-A3E3-723BEA898919}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">Communication Matrices</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">70</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{A722E2B8-21FF-45CB-86EB-A3414D49D7AF}</EntityID>
			<Targets/>
		</item>
		<item>
			<DisplayName type="key">External Cable Harness</DisplayName>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">131328</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">32</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{8ABE8996-5BA4-4722-B7A8-BDFE8EEE5CEC}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Application.cfgx</Name>
			<DisplayName type="key">Core Application</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">260</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">20</Type>
			<ItemInfoDate type="key">28.03.2024 10:08:15</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{84666013-649B-4E59-93A0-9A9A085B0984}</EntityID>
			<Targets/>
		</item>
		<item>
			<Name type="key">Build Results</Name>
			<DisplayName type="key">Build Results</DisplayName>
			<Path type="key">.</Path>
			<Component type="key">ProjectApplication</Component>
			<Flags type="key">256</Flags>
			<ExtendedFlags type="key">0</ExtendedFlags>
			<Type type="key">58</Type>
			<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
			<ItemInfoPath type="key"/>
			<ItemInfoDocs type="key"/>
			<ItemInfoDescr type="key"/>
			<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
			<ItemInfoAddInfoDb type="key"/>
			<Log type="key"/>
			<DatabaseID type="key">-1</DatabaseID>
			<EntityID type="key">{725495FA-E03C-4E55-998B-21915B393C59}</EntityID>
			<Targets/>
			<item>
				<Name type="key">Build Results</Name>
				<DisplayName type="key">itSDFROOT</DisplayName>
				<Path type="key">.</Path>
				<Component type="key">ProjectApplication</Component>
				<Flags type="key">260</Flags>
				<ExtendedFlags type="key">0</ExtendedFlags>
				<Type type="key">29</Type>
				<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
				<ItemInfoPath type="key"/>
				<ItemInfoDocs type="key"/>
				<ItemInfoDescr type="key"/>
				<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
				<ItemInfoAddInfoDb type="key"/>
				<Log type="key"/>
				<DatabaseID type="key">-1</DatabaseID>
				<EntityID type="key">{F6B6BAC5-EB44-4285-BEDC-EC5BD2870091}</EntityID>
				<Targets/>
				<item>
					<Name type="key">Furuta_Acados.dsbuildinfo</Name>
					<DisplayName type="key">Furuta_Acados.dsbuildinfo</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">260</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">4</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{8E3761E0-460B-4AE1-A22C-6657E2D8A000}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Furuta_Acados.rta</Name>
					<DisplayName type="key">Furuta_Acados.rta</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">37</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{15F3E3FE-1655-4E5F-8F53-AEBE674F9A76}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Furuta_Acados.sdf</Name>
					<DisplayName type="key">Furuta_Acados.sdf</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">35</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{4B15C3A1-AB00-44B3-87F3-6167842EB54B}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Furuta_Model.expswcfg</Name>
					<DisplayName type="key">Furuta_Model.expswcfg</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">71</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{2A7198B5-F45C-4972-9378-19DD610B00D7}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Furuta_Model.map</Name>
					<DisplayName type="key">Furuta_Model.map</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">36</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{A7538352-8737-42D4-84E5-1CFC7C83B3D8}</EntityID>
					<Targets/>
				</item>
				<item>
					<Name type="key">Furuta_Model.trc</Name>
					<DisplayName type="key">Furuta_Model.trc</DisplayName>
					<Path type="key">.\Build Results</Path>
					<Component type="key">ProjectApplication</Component>
					<Flags type="key">256</Flags>
					<ExtendedFlags type="key">0</ExtendedFlags>
					<Type type="key">34</Type>
					<ItemInfoDate type="key">28.03.2024 10:29:47</ItemInfoDate>
					<ItemInfoPath type="key"/>
					<ItemInfoDocs type="key"/>
					<ItemInfoDescr type="key"/>
					<ItemInfoAuthor type="key">Administrator</ItemInfoAuthor>
					<ItemInfoAddInfoDb type="key"/>
					<Log type="key"/>
					<DatabaseID type="key">-1</DatabaseID>
					<EntityID type="key">{4C7B9F3D-B3FB-4A95-8A24-458F3C6CA88D}</EntityID>
					<Targets/>
				</item>
			</item>
		</item>
	</application>
</Root>